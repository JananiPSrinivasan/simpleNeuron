module mac(
    input logic signed [7:0] x,
    input logic signed [7:0] weight,
    output logic signed [7:0]
);
endmodule